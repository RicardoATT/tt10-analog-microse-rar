magic
tech sky130A
magscale 1 2
timestamp 1740782616
<< error_p >>
rect -29 123 29 129
rect -29 89 -17 123
rect -29 83 29 89
rect -67 24 -21 36
rect -67 -24 -61 24
rect -67 -36 -21 -24
rect -29 -89 29 -83
rect -29 -123 -17 -89
rect -29 -129 29 -123
<< nwell >>
rect -211 -261 211 261
<< pmoshvt >>
rect -15 -42 15 42
<< pdiff >>
rect -73 30 -15 42
rect -73 -30 -61 30
rect -27 -30 -15 30
rect -73 -42 -15 -30
rect 15 30 73 42
rect 15 -30 27 30
rect 61 -30 73 30
rect 15 -42 73 -30
<< pdiffc >>
rect -61 -30 -27 30
rect 27 -30 61 30
<< nsubdiff >>
rect -175 191 175 225
rect -175 -191 -141 191
rect 141 -191 175 191
rect -175 -225 -79 -191
rect 79 -225 175 -191
<< nsubdiffcont >>
rect -79 -225 79 -191
<< poly >>
rect -33 123 33 139
rect -33 89 -17 123
rect 17 89 33 123
rect -33 73 33 89
rect -15 42 15 73
rect -15 -73 15 -42
rect -33 -89 33 -73
rect -33 -123 -17 -89
rect 17 -123 33 -89
rect -33 -139 33 -123
<< polycont >>
rect -17 89 17 123
rect -17 -123 17 -89
<< locali >>
rect -33 89 -17 123
rect 17 89 33 123
rect -61 30 -27 46
rect -61 -46 -27 -30
rect 27 30 61 46
rect 27 -46 61 -30
rect -33 -123 -17 -89
rect 17 -123 33 -89
rect -95 -225 -79 -191
rect 79 -225 95 -191
<< viali >>
rect -17 89 17 123
rect -61 -24 -27 24
rect 27 -30 61 30
rect -17 -123 17 -89
<< metal1 >>
rect -29 123 29 129
rect -29 89 -17 123
rect 17 89 29 123
rect -29 83 29 89
rect -67 24 -21 36
rect -67 -24 -61 24
rect -27 -24 -21 24
rect -67 -36 -21 -24
rect 21 30 67 42
rect 21 -30 27 30
rect 61 -30 67 30
rect 21 -42 67 -30
rect -29 -89 29 -83
rect -29 -123 -17 -89
rect 17 -123 29 -89
rect -29 -129 29 -123
<< properties >>
string FIXED_BBOX -158 -208 158 208
string gencell sky130_fd_pr__pfet_01v8_hvt
string library sky130
string parameters w 0.42 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 80 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
