magic
tech sky130A
magscale 1 2
timestamp 1740881680
<< nwell >>
rect 1930 176 1986 242
rect 2144 -25 2178 257
<< pwell >>
rect 1068 177 1237 243
rect 1915 -949 2286 -893
<< locali >>
rect 2144 473 2197 512
rect 1136 349 2157 383
rect 1622 294 1656 349
rect 1099 -126 1133 124
rect 1622 69 1656 127
rect 1622 35 1832 69
rect 1622 -38 1656 35
rect 2144 -25 2178 257
rect 1622 -72 1832 -38
rect 1622 -122 1656 -72
rect 1099 -352 1134 -300
rect 1301 -352 1336 -350
rect 1099 -387 1336 -352
rect 1099 -971 1134 -387
rect 1348 -510 1550 -485
rect 1622 -510 1656 -298
rect 1348 -519 1656 -510
rect 1516 -550 1656 -519
rect 2144 -969 2178 -724
rect 1108 -1152 1124 -1136
rect 1100 -1178 1134 -1152
rect 1604 -1178 1638 -1136
rect 2144 -1178 2178 -1144
rect 1027 -1187 2398 -1178
rect 1061 -1212 2398 -1187
<< viali >>
rect 2197 473 2236 512
rect 1102 349 1136 383
rect 1832 35 1866 69
rect 1832 -72 1866 -38
rect 1301 -350 1336 -315
rect 1314 -519 1348 -485
rect 1027 -1221 1061 -1187
rect 2398 -1212 2432 -1178
<< metal1 >>
rect 2191 512 2242 524
rect 2191 473 2197 512
rect 2236 485 2281 512
rect 2476 500 2785 533
rect 2236 479 2288 485
rect 2191 461 2236 473
rect 2476 473 2509 500
rect 2236 421 2288 427
rect 2568 438 2624 446
rect 1096 383 1142 395
rect 1033 349 1102 383
rect 1136 349 1142 383
rect 2400 391 2452 397
rect 1823 367 2286 370
rect 1096 337 1142 349
rect 1291 319 2286 367
rect 2568 382 2654 438
rect 2710 382 2716 438
rect 2568 380 2624 382
rect 2400 333 2452 339
rect 1291 277 1339 319
rect 1285 271 1345 277
rect 1068 177 1242 243
rect 1279 237 1351 271
rect 1186 122 1242 177
rect 1180 66 1186 122
rect 1242 66 1248 122
rect 1185 -195 1241 -179
rect 1283 -185 1355 183
rect 1389 177 1445 243
rect 1724 242 1761 319
rect 1708 176 1764 242
rect 1823 236 1871 319
rect 2230 251 2286 319
rect 2752 292 2785 500
rect 1832 75 1866 182
rect 1930 176 1986 242
rect 2230 189 2286 195
rect 1820 69 1878 75
rect 1820 35 1832 69
rect 1866 35 1878 69
rect 1820 29 1878 35
rect 2345 31 2386 292
rect 2498 246 2785 292
rect 2238 -6 2386 31
rect 2233 -10 2386 -6
rect 2233 -12 2285 -10
rect 1826 -38 1872 -26
rect 1816 -72 1832 -38
rect 1866 -72 1878 -38
rect 2233 -70 2285 -64
rect 2472 -35 2796 2
rect 2472 -65 2509 -35
rect 1035 -229 1241 -195
rect 1185 -245 1241 -229
rect 1301 -240 1336 -239
rect 1288 -315 1348 -240
rect 1389 -245 1445 -179
rect 1708 -246 1764 -180
rect 1816 -182 1878 -72
rect 2568 -85 2624 -80
rect 2380 -134 2432 -128
rect 1288 -350 1301 -315
rect 1336 -350 1348 -315
rect 1289 -356 1348 -350
rect 1723 -406 1758 -246
rect 1034 -441 1758 -406
rect 1308 -485 1354 -473
rect 1186 -514 1242 -508
rect 1308 -519 1314 -485
rect 1348 -519 1354 -485
rect 1308 -531 1354 -519
rect 1094 -740 1150 -734
rect 1027 -796 1094 -740
rect 1094 -802 1150 -796
rect 1186 -1090 1242 -570
rect 1314 -604 1348 -531
rect 1289 -828 1358 -662
rect 1408 -670 1464 -604
rect 1594 -669 1774 -600
rect 1811 -608 1877 -240
rect 1930 -246 1986 -180
rect 2230 -303 2286 -176
rect 2432 -180 2464 -139
rect 2568 -141 2665 -85
rect 2721 -141 2727 -85
rect 2568 -146 2624 -141
rect 2380 -192 2432 -186
rect 2759 -234 2796 -35
rect 2282 -355 2286 -303
rect 1594 -828 1663 -669
rect 1289 -897 1663 -828
rect 1811 -893 1873 -662
rect 1930 -668 1986 -602
rect 2230 -740 2286 -355
rect 2394 -592 2455 -253
rect 2502 -266 2796 -234
rect 2502 -280 2795 -266
rect 2230 -802 2286 -796
rect 1289 -1030 1358 -897
rect 1784 -949 2286 -893
rect 1286 -1172 1346 -1084
rect 1390 -1090 1446 -1024
rect 1690 -1090 1746 -1024
rect 1784 -1030 1844 -949
rect 1894 -1090 1950 -949
rect 2230 -1089 2286 -949
rect 2389 -1021 2454 -666
rect 2550 -668 2606 -602
rect 1790 -1172 1850 -1092
rect 2398 -1166 2432 -1089
rect 2550 -1090 2606 -1024
rect 998 -1187 1850 -1172
rect 998 -1221 1027 -1187
rect 1061 -1221 1850 -1187
rect 998 -1232 1850 -1221
rect 2392 -1178 2438 -1166
rect 2392 -1212 2398 -1178
rect 2432 -1212 2438 -1178
rect 2392 -1224 2438 -1212
rect 1021 -1233 1067 -1232
<< via1 >>
rect 2236 427 2288 479
rect 2400 339 2452 391
rect 2654 382 2710 438
rect 1186 66 1242 122
rect 2230 195 2286 251
rect 2233 -64 2285 -12
rect 1186 -570 1242 -514
rect 1094 -796 1150 -740
rect 2380 -186 2432 -134
rect 2665 -141 2721 -85
rect 2230 -355 2282 -303
rect 2230 -796 2286 -740
<< metal2 >>
rect 2230 427 2236 479
rect 2288 427 2294 479
rect 2654 438 2710 444
rect 2243 384 2282 427
rect 2394 384 2400 391
rect 2243 345 2400 384
rect 2394 339 2400 345
rect 2452 339 2458 391
rect 2224 195 2230 251
rect 2286 209 2292 251
rect 2654 209 2710 382
rect 2286 195 2710 209
rect 2230 153 2710 195
rect 1186 122 1242 128
rect 1186 -514 1242 66
rect 2227 -64 2233 -12
rect 2285 -64 2291 -12
rect 2239 -140 2280 -64
rect 2665 -85 2721 -79
rect 2374 -140 2380 -134
rect 2239 -181 2380 -140
rect 2374 -186 2380 -181
rect 2432 -186 2438 -134
rect 2665 -147 2721 -141
rect 2667 -303 2719 -147
rect 2224 -355 2230 -303
rect 2282 -355 2719 -303
rect 1180 -570 1186 -514
rect 1242 -570 1248 -514
rect 1088 -796 1094 -740
rect 1150 -796 2230 -740
rect 2286 -796 2292 -740
use sky130_fd_pr__nfet_01v8_LAQ5H5  XM7
timestamp 1740782616
transform 0 1 2418 1 0 -635
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_LY9833  XM8
timestamp 1740782616
transform 0 1 1315 1 0 -212
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_JC5RM4  XM9
timestamp 1740782616
transform 0 1 2427 1 0 -161
box -263 -319 263 319
use sky130_fd_pr__pfet_01v8_JC5RM4  XM10
timestamp 1740782616
transform 0 1 2427 1 0 365
box -263 -319 263 319
use sky130_fd_pr__pfet_01v8_EBBUFJ  XM11
timestamp 1740782616
transform 0 -1 1325 1 0 -635
box -211 -261 211 261
use sky130_fd_pr__nfet_01v8_LY9833  XM12
timestamp 1740782616
transform 0 1 1316 1 0 -1057
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_hvt_EBBUFJ  XM13
timestamp 1740782616
transform 0 1 1847 1 0 -635
box -211 -261 211 261
use sky130_fd_pr__nfet_01v8_lvt_LAQ5H5
timestamp 1740782616
transform 0 1 2418 1 0 -1057
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_LY9833  XM16
timestamp 1740782616
transform 0 1 1820 1 0 -1057
box -211 -252 211 252
use sky130_fd_pr__pfet_01v8_hvt_EBBUFJ  XM17
timestamp 1740782616
transform 0 1 1847 -1 0 209
box -211 -261 211 261
use sky130_fd_pr__pfet_01v8_EBBUFJ  XM18
timestamp 1740782616
transform 0 1 1847 1 0 -213
box -211 -261 211 261
use sky130_fd_pr__nfet_01v8_lvt_LY9833  XM19
timestamp 1740782616
transform 0 1 1315 1 0 210
box -211 -252 211 252
<< labels >>
flabel metal1 s 1049 365 1049 365 0 FreeSans 240 0 0 0 vdd
port 5 nsew
flabel metal1 s 1049 -214 1049 -214 0 FreeSans 240 0 0 0 exc_ctrl
port 4 nsew
flabel locali s 1043 -425 1043 -425 0 FreeSans 240 0 0 0 inh_ctrl
port 3 nsew
flabel metal1 1214 -867 1216 -864 0 FreeSans 240 0 0 0 input_syn
port 2 nsew
flabel metal1 1014 -1201 1014 -1201 0 FreeSans 240 0 0 0 GND
port 1 nsew
flabel metal1 s 1047 -768 1047 -768 0 FreeSans 240 0 0 0 syps_ctrl
port 6 nsew
flabel metal1 s 2426 -434 2426 -434 0 FreeSans 240 0 0 0 output_syps
port 7 nsew
<< end >>
