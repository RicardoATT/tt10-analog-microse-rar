magic
tech sky130A
magscale 1 2
timestamp 1740946172
<< metal1 >>
rect 4353 41687 4359 41739
rect 4411 41729 4417 41739
rect 4411 41696 4929 41729
rect 4411 41687 4417 41696
rect 4751 41695 4929 41696
rect 4676 41654 4732 41660
rect 4676 40606 4732 41598
rect 4827 41523 4833 41589
rect 4899 41523 4996 41589
rect 4786 41108 4792 41160
rect 4844 41151 4850 41160
rect 4844 41117 4931 41151
rect 4844 41108 4850 41117
rect 4871 40905 4931 40940
rect 4871 40837 4906 40905
rect 6256 40876 6686 40937
rect 4863 40831 4915 40837
rect 4863 40773 4915 40779
rect 4676 40550 4945 40606
rect 4211 40112 4217 40170
rect 4275 40112 4903 40170
rect 6625 40061 6686 40876
rect 4560 40000 6686 40061
rect 4560 2179 4621 40000
rect 4560 2118 18840 2179
rect 18779 1829 18840 2118
rect 18779 1762 18840 1768
<< via1 >>
rect 4359 41687 4411 41739
rect 4676 41598 4732 41654
rect 4833 41523 4899 41589
rect 4792 41108 4844 41160
rect 4863 40779 4915 40831
rect 4217 40112 4275 40170
rect 18779 1768 18840 1829
<< metal2 >>
rect 27449 44362 27458 44364
rect 4676 44306 27458 44362
rect 2266 41684 2275 41744
rect 2335 41730 2344 41744
rect 4359 41739 4411 41745
rect 2335 41697 4359 41730
rect 2335 41684 2344 41697
rect 4359 41681 4411 41687
rect 4676 41654 4732 44306
rect 27449 44304 27458 44306
rect 27518 44304 27527 44364
rect 4670 41598 4676 41654
rect 4732 41598 4738 41654
rect 4833 41589 4899 41595
rect 4833 41511 4899 41523
rect 4553 41445 4899 41511
rect 2165 40111 2174 40171
rect 2234 40170 2243 40171
rect 4217 40170 4275 40176
rect 2234 40112 4217 40170
rect 2234 40111 2243 40112
rect 4217 40106 4275 40112
rect 4553 2183 4619 41445
rect 4792 41160 4844 41166
rect 4701 41117 4792 41151
rect 4701 2309 4735 41117
rect 4792 41102 4844 41108
rect 4857 40779 4863 40831
rect 4915 40779 4921 40831
rect 4872 2412 4907 40779
rect 4872 2377 30455 2412
rect 4701 2275 26619 2309
rect 4553 2117 22745 2183
rect 18773 1768 18779 1829
rect 18840 1768 18846 1829
rect 18779 1373 18840 1768
rect 22679 1731 22745 2117
rect 26585 2009 26619 2275
rect 30420 2084 30455 2377
rect 30408 2075 30468 2084
rect 26572 2000 26632 2009
rect 30408 2006 30468 2015
rect 26572 1931 26632 1940
rect 22679 1656 22745 1665
rect 18779 1303 18840 1312
<< via2 >>
rect 2275 41684 2335 41744
rect 27458 44304 27518 44364
rect 2174 40111 2234 40171
rect 30408 2015 30468 2075
rect 26572 1940 26632 2000
rect 22679 1665 22745 1731
rect 18779 1312 18840 1373
<< metal3 >>
rect 27654 44692 27660 44756
rect 27724 44692 27730 44756
rect 27453 44364 27523 44369
rect 27662 44364 27722 44692
rect 27453 44304 27458 44364
rect 27518 44304 27722 44364
rect 27453 44299 27523 44304
rect 354 41682 360 41746
rect 424 41744 430 41746
rect 2270 41744 2340 41749
rect 424 41684 2275 41744
rect 2335 41684 2340 41744
rect 424 41682 430 41684
rect 2270 41679 2340 41684
rect 1808 40109 1814 40173
rect 1878 40171 1884 40173
rect 2169 40171 2239 40176
rect 1878 40111 2174 40171
rect 2234 40111 2239 40171
rect 1878 40109 1884 40111
rect 2169 40106 2239 40111
rect 30403 2075 30473 2080
rect 30403 2015 30408 2075
rect 30468 2015 30473 2075
rect 30403 2010 30473 2015
rect 26567 2000 26637 2005
rect 26567 1940 26572 2000
rect 26632 1940 26637 2000
rect 26567 1935 26637 1940
rect 22674 1731 22750 1736
rect 22674 1665 22679 1731
rect 22745 1665 22750 1731
rect 22674 1660 22750 1665
rect 18774 1373 18845 1378
rect 18774 1312 18779 1373
rect 18840 1312 18845 1373
rect 18774 1307 18845 1312
rect 18779 613 18840 1307
rect 22679 841 22745 1660
rect 22679 769 22745 775
rect 26572 686 26632 1935
rect 30408 1090 30468 2010
rect 30406 1084 30470 1090
rect 30406 1014 30470 1020
rect 26570 680 26634 686
rect 18778 607 18842 613
rect 26570 610 26634 616
rect 18778 537 18842 543
<< via3 >>
rect 27660 44692 27724 44756
rect 360 41682 424 41746
rect 1814 40109 1878 40173
rect 22679 775 22745 841
rect 30406 1020 30470 1084
rect 26570 616 26634 680
rect 18778 543 18842 607
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44757 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 27659 44756 27725 44757
rect 27659 44692 27660 44756
rect 27724 44692 27725 44756
rect 27659 44691 27725 44692
rect 200 41746 600 44152
rect 200 41682 360 41746
rect 424 41682 600 41746
rect 200 1000 600 41682
rect 800 40171 1200 44152
rect 1813 40173 1879 40174
rect 1813 40171 1814 40173
rect 800 40111 1814 40171
rect 800 1000 1200 40111
rect 1813 40109 1814 40111
rect 1878 40109 1879 40173
rect 1813 40108 1879 40109
rect 30405 1084 30471 1085
rect 30405 1020 30406 1084
rect 30470 1020 30471 1084
rect 30405 1019 30471 1020
rect 22678 841 22746 842
rect 22678 775 22679 841
rect 22745 775 22746 841
rect 22678 774 22746 775
rect 18777 607 18843 608
rect 18777 543 18778 607
rect 18842 543 18843 607
rect 18777 542 18843 543
rect 18780 200 18841 542
rect 22679 200 22745 774
rect 26569 680 26635 681
rect 26569 616 26570 680
rect 26634 616 26635 680
rect 26569 615 26635 616
rect 26572 200 26632 615
rect 30408 200 30468 1019
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 200
use synapse  synapse_0
timestamp 1740881680
transform 1 0 3862 0 1 41346
box 998 -1268 2796 628
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
